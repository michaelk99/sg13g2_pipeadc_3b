.save @n.xamp1.xmn1.nsg13_lv_nmos[ids]
.save @n.xamp1.xmn1.nsg13_lv_nmos[vth]
.save @n.xamp1.xmn1.nsg13_lv_nmos[vgs]
.save @n.xamp1.xmn1.nsg13_lv_nmos[vds]
.save @n.xamp1.xmn1.nsg13_lv_nmos[vdss]
.save @n.xamp1.xmn1.nsg13_lv_nmos[gm]
.save @n.xamp1.xmn1.nsg13_lv_nmos[gds]
.save @n.xamp1.xmn1.nsg13_lv_nmos[cgs]
.save @n.xamp1.xmn1.nsg13_lv_nmos[cgg]

.save @n.xamp1.xmn2.nsg13_lv_nmos[ids]
.save @n.xamp1.xmn2.nsg13_lv_nmos[vth]
.save @n.xamp1.xmn2.nsg13_lv_nmos[vgs]
.save @n.xamp1.xmn2.nsg13_lv_nmos[vds]
.save @n.xamp1.xmn2.nsg13_lv_nmos[vdss]
.save @n.xamp1.xmn2.nsg13_lv_nmos[gm]
.save @n.xamp1.xmn2.nsg13_lv_nmos[gds]
.save @n.xamp1.xmn2.nsg13_lv_nmos[cgs]
.save @n.xamp1.xmn2.nsg13_lv_nmos[cgg]

.save @n.xamp1.xmn3.nsg13_lv_nmos[ids]
.save @n.xamp1.xmn3.nsg13_lv_nmos[vth]
.save @n.xamp1.xmn3.nsg13_lv_nmos[vgs]
.save @n.xamp1.xmn3.nsg13_lv_nmos[vds]
.save @n.xamp1.xmn3.nsg13_lv_nmos[vdss]
.save @n.xamp1.xmn3.nsg13_lv_nmos[gm]
.save @n.xamp1.xmn3.nsg13_lv_nmos[gds]
.save @n.xamp1.xmn3.nsg13_lv_nmos[cgs]
.save @n.xamp1.xmn3.nsg13_lv_nmos[cgg]

.save @n.xamp1.xmn4.nsg13_lv_nmos[ids]
.save @n.xamp1.xmn4.nsg13_lv_nmos[vth]
.save @n.xamp1.xmn4.nsg13_lv_nmos[vgs]
.save @n.xamp1.xmn4.nsg13_lv_nmos[vds]
.save @n.xamp1.xmn4.nsg13_lv_nmos[vdss]
.save @n.xamp1.xmn4.nsg13_lv_nmos[gm]
.save @n.xamp1.xmn4.nsg13_lv_nmos[gds]
.save @n.xamp1.xmn4.nsg13_lv_nmos[cgs]
.save @n.xamp1.xmn4.nsg13_lv_nmos[cgg]







.save @n.xamp1.xmp1.nsg13_lv_pmos[ids]
.save @n.xamp1.xmp1.nsg13_lv_pmos[vth]
.save @n.xamp1.xmp1.nsg13_lv_pmos[vgs]
.save @n.xamp1.xmp1.nsg13_lv_pmos[vds]
.save @n.xamp1.xmp1.nsg13_lv_pmos[vdss]
.save @n.xamp1.xmp1.nsg13_lv_pmos[gm]
.save @n.xamp1.xmp1.nsg13_lv_pmos[gds]
.save @n.xamp1.xmp1.nsg13_lv_pmos[cgs]
.save @n.xamp1.xmp1.nsg13_lv_pmos[cgg]

.save @n.xamp1.xmp2.nsg13_lv_pmos[ids]
.save @n.xamp1.xmp2.nsg13_lv_pmos[vth]
.save @n.xamp1.xmp2.nsg13_lv_pmos[vgs]
.save @n.xamp1.xmp2.nsg13_lv_pmos[vds]
.save @n.xamp1.xmp2.nsg13_lv_pmos[vdss]
.save @n.xamp1.xmp2.nsg13_lv_pmos[gm]
.save @n.xamp1.xmp2.nsg13_lv_pmos[gds]
.save @n.xamp1.xmp2.nsg13_lv_pmos[cgs]
.save @n.xamp1.xmp2.nsg13_lv_pmos[cgg]

.save @n.xamp1.xmp3.nsg13_lv_pmos[ids]
.save @n.xamp1.xmp3.nsg13_lv_pmos[vth]
.save @n.xamp1.xmp3.nsg13_lv_pmos[vgs]
.save @n.xamp1.xmp3.nsg13_lv_pmos[vds]
.save @n.xamp1.xmp3.nsg13_lv_pmos[vdss]
.save @n.xamp1.xmp3.nsg13_lv_pmos[gm]
.save @n.xamp1.xmp3.nsg13_lv_pmos[gds]
.save @n.xamp1.xmp3.nsg13_lv_pmos[cgs]
.save @n.xamp1.xmp3.nsg13_lv_pmos[cgg]
